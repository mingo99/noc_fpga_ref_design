//////////////////////////////////////
// ACE GENERATED VERILOG INCLUDE FILE
// Generated on: 2021.05.04 at 06:44:45 PDT
// By: ACE 8.3.3
// From project: pcie_ref_design_top
//////////////////////////////////////
// User Design Signal List Include File
//////////////////////////////////////

    // Ports for clock_io_bank
    // Ports for gpio_bank_north
    logic        i_reset_n;
    logic        i_start;
    logic        o_fail;
    logic        o_fail_oe;
    logic        o_mstr_test_complete;
    logic        o_mstr_test_complete_oe;
    // Ports for noc
    // Ports for pci_express_x16
    // Status
    logic  [3:0] pci_express_x16_status_flr_pf_active;
    logic        pci_express_x16_status_flr_vf_active;
    logic  [5:0] pci_express_x16_status_ltssm_state;
    // Ports for pci_express_x8
    // Status
    logic  [5:0] pci_express_x8_status_ltssm_state;
    // Ports for pll_1
    logic        i_clk;
    logic        pll_1_lock;

//////////////////////////////////////
// End User Design Signal List Include File
//////////////////////////////////////
