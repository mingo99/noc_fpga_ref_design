//////////////////////////////////////
// ACE GENERATED VERILOG INCLUDE FILE
// Generated on: 2022.01.10 at 23:18:52 PST
// By: ACE 8.6.1
// From project: noc_2d_ref_design_top
//////////////////////////////////////
// User Design Port List Include File
//////////////////////////////////////

    // Ports for noc_2d
    // Ports for pll_chk_clk
    input        i_chk_clk,
    input        pll_chk_clk_lock,
    // Ports for pll_send_clk
    input        i_cc_clk,
    input        i_reg_clk,
    input        i_send_clk,
    input        pll_send_clk_lock,
    // Ports for vp_1550_clkio_ne
    input        fpga_rst_l,
    // Ports for vp_1550_clkio_nw
    // Ports for vp_1550_clkio_se
    // Ports for vp_1550_clkio_sw
    // Ports for vp_1550_gpio_n_b0
    input        ext_gpio_fpga_in[0],
    input        ext_gpio_fpga_in[1],
    input        ext_gpio_fpga_in[2],
    input        ext_gpio_fpga_in[3],
    input        ext_gpio_fpga_in[4],
    input        ext_gpio_fpga_in[5],
    input        ext_gpio_fpga_in[6],
    input        ext_gpio_fpga_in[7],
    output       ext_gpio_fpga_oe[0],
    output       ext_gpio_fpga_oe[1],
    output       ext_gpio_fpga_oe[2],
    output       ext_gpio_fpga_oe[3],
    output       ext_gpio_fpga_oe[4],
    output       ext_gpio_fpga_oe[5],
    output       ext_gpio_fpga_oe[6],
    output       ext_gpio_fpga_oe[7],
    output       ext_gpio_fpga_out[0],
    output       ext_gpio_fpga_out[1],
    output       ext_gpio_fpga_out[2],
    output       ext_gpio_fpga_out[3],
    output       ext_gpio_fpga_out[4],
    output       ext_gpio_fpga_out[5],
    output       ext_gpio_fpga_out[6],
    output       ext_gpio_fpga_out[7],
    output       ext_gpio_oe_l,
    output       ext_gpio_oe_l_oe,
    output       led_oe_l,
    output       led_oe_l_oe,
    // Ports for vp_1550_gpio_n_b1
    output       ext_gpio_dir[0],
    output       ext_gpio_dir[1],
    output       ext_gpio_dir[2],
    output       ext_gpio_dir[3],
    output       ext_gpio_dir[4],
    output       ext_gpio_dir[5],
    output       ext_gpio_dir[6],
    output       ext_gpio_dir[7],
    output       ext_gpio_dir_oe[0],
    output       ext_gpio_dir_oe[1],
    output       ext_gpio_dir_oe[2],
    output       ext_gpio_dir_oe[3],
    output       ext_gpio_dir_oe[4],
    output       ext_gpio_dir_oe[5],
    output       ext_gpio_dir_oe[6],
    output       ext_gpio_dir_oe[7],
    output       led_l[4],
    output       led_l[5],
    output       led_l_oe[4],
    output       led_l_oe[5],
    // Ports for vp_1550_gpio_n_b2
    output       led_l[0],
    output       led_l[1],
    output       led_l[2],
    output       led_l[3],
    output       led_l[6],
    output       led_l[7],
    output       led_l_oe[0],
    output       led_l_oe[1],
    output       led_l_oe[2],
    output       led_l_oe[3],
    output       led_l_oe[6],
    output       led_l_oe[7],
    // Ports for vp_1550_gpio_s_b0
    input        fpga_avr_rxd,
    input        fpga_ftdi_rxd,
    input        fpga_i2c_mux_gnt,
    input        irq_to_fpga,
    input        qsfp_int_fpga_l,
    output       fpga_avr_txd,
    output       fpga_avr_txd_oe,
    output       fpga_ftdi_txd,
    output       fpga_ftdi_txd_oe,
    output       fpga_i2c_req_l,
    output       fpga_i2c_req_l_oe,
    output       irq_to_avr,
    output       irq_to_avr_oe,
    output       test[1],
    output       test_oe[1],
    // Ports for vp_1550_gpio_s_b1
    input        mcio_vio_45_10_clk,
    input        mcio_vio_in[0],
    input        mcio_vio_in[1],
    input        mcio_vio_in[2],
    input        mcio_vio_in[3],
    output       mcio_dir[0],
    output       mcio_dir[1],
    output       mcio_dir[2],
    output       mcio_dir[3],
    output       mcio_dir_45,
    output       mcio_dir_45_oe,
    output       mcio_dir_oe[0],
    output       mcio_dir_oe[1],
    output       mcio_dir_oe[2],
    output       mcio_dir_oe[3],
    output       mcio_vio_oe[0],
    output       mcio_vio_oe[1],
    output       mcio_vio_oe[2],
    output       mcio_vio_oe[3],
    output       mcio_vio_out[0],
    output       mcio_vio_out[1],
    output       mcio_vio_out[2],
    output       mcio_vio_out[3],
    output       test[2],
    output       test_oe[2],
    // Ports for vp_1550_gpio_s_b2
    input        fpga_sys_scl_in,
    input        fpga_sys_sda_in,
    input        mcio_scl_in,
    input        mcio_sda_in,
    output       fpga_sys_scl_oe,
    output       fpga_sys_scl_out,
    output       fpga_sys_sda_oe,
    output       fpga_sys_sda_out,
    output       mcio_oe1_l,
    output       mcio_oe1_l_oe,
    output       mcio_oe_45_l,
    output       mcio_oe_45_l_oe,
    output       mcio_scl_oe,
    output       mcio_scl_out,
    output       mcio_sda_oe,
    output       mcio_sda_out,
    // Ports for vp_1550_pll_nw_2
    input        pll_nw_2_ref0_312p5_clk,
    input        vp_1550_pll_nw_2_lock,
    // Ports for vp_1550_pll_sw_2
    input        pll_sw_2_ref1_312p5_clk,
    input        vp_1550_pll_sw_2_lock 

//////////////////////////////////////
// End User Design Port List Include File
//////////////////////////////////////
