// Include before other files, to turn off the default nettype. This enforces
// use of proper declarations (recommended).

`default_nettype none
